-- Copyright of the original ROM contents respectfully acknowleged

-- This file was created and maintaned by Grant Searle 2014
-- You are free to use this file in your own projects but must never charge for it nor use it without
-- acknowledgement.
-- Please ask permission from Grant Searle before republishing elsewhere.
-- If you use this file or any part of it, please add an acknowledgement to myself and
-- a link back to my main web site http://searle.hostei.com/grant/    
-- and to the UK101 page at http://searle.hostei.com/grant/uk101FPGA/index.html
--
-- Please check on the above web pages to see if there are any updates before using this file.
-- If for some reason the page is no longer available, please search for "Grant Searle"
-- on the internet to see if I have moved to another web hosting service.
--
-- Grant Searle
-- eMail address available on my main web page link above.


library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	use ieee.std_logic_unsigned.all;

ENTITY CegmonRom IS

	PORT
	(
		address : in std_logic_vector(10 downto 0);
		q : out std_logic_vector(7 downto 0)
	);
END CegmonRom;

architecture behavior of CegmonRom is
type romtable is array (0 to 2047) of std_logic_vector(7 downto 0);
constant romdata : romtable :=
(
x"86",x"30",x"84",x"31",x"85",x"34",x"A5",x"34",
x"30",x"42",x"A5",x"31",x"85",x"37",x"A5",x"30",
x"85",x"36",x"86",x"3E",x"A5",x"30",x"85",x"32",
x"29",x"07",x"AA",x"A5",x"31",x"49",x"FF",x"4A",
x"66",x"32",x"4A",x"66",x"32",x"4A",x"66",x"32",
x"09",x"80",x"85",x"33",x"A5",x"34",x"4A",x"BD",
x"43",x"F8",x"A2",x"00",x"90",x"04",x"01",x"32",
x"D0",x"04",x"49",x"FF",x"21",x"32",x"81",x"32",
x"A6",x"3E",x"60",x"80",x"40",x"20",x"10",x"08",
x"04",x"02",x"01",x"00",x"A2",x"02",x"B5",x"2F",
x"EA",x"38",x"F5",x"35",x"B0",x"05",x"49",x"FF",
x"69",x"01",x"18",x"95",x"37",x"66",x"35",x"CA",
x"D0",x"EC",x"A5",x"38",x"D0",x"04",x"C5",x"39",
x"F0",x"0B",x"0A",x"B0",x"07",x"06",x"39",x"90",
x"F9",x"66",x"39",x"18",x"6A",x"85",x"38",x"A0",
x"00",x"A2",x"00",x"8A",x"38",x"65",x"38",x"AA",
x"90",x"0A",x"24",x"35",x"30",x"04",x"E6",x"30",
x"D0",x"02",x"C6",x"30",x"98",x"38",x"65",x"39",
x"A8",x"90",x"0A",x"24",x"35",x"70",x"04",x"E6",
x"31",x"D0",x"02",x"C6",x"31",x"20",x"12",x"F8",
x"A5",x"30",x"C5",x"36",x"D0",x"D5",x"A5",x"31",
x"C5",x"37",x"D0",x"CF",x"60",x"A9",x"40",x"85",
x"E0",x"A9",x"D0",x"85",x"E1",x"A9",x"03",x"8D",
x"00",x"F0",x"A9",x"11",x"4C",x"96",x"FB",x"60",
x"48",x"AD",x"00",x"F0",x"4A",x"4A",x"90",x"F9",
x"68",x"8D",x"01",x"F0",x"60",x"49",x"FF",x"8D",
x"00",x"DF",x"49",x"FF",x"60",x"48",x"20",x"DE",
x"F8",x"AA",x"68",x"CA",x"E8",x"60",x"AD",x"00",
x"DF",x"49",x"FF",x"60",x"A2",x"02",x"BD",x"DB",
x"FF",x"95",x"BC",x"CA",x"10",x"F8",x"4C",x"00",
x"00",x"A0",x"09",x"B9",x"AC",x"FC",x"99",x"06",
x"02",x"88",x"D0",x"F7",x"A2",x"04",x"4C",x"07",
x"02",x"C8",x"D0",x"FA",x"EE",x"09",x"02",x"EE",
x"0C",x"02",x"CA",x"D0",x"F1",x"A0",x"1F",x"A9",
x"60",x"99",x"E0",x"D3",x"88",x"10",x"FA",x"60",
x"68",x"85",x"E2",x"68",x"68",x"68",x"68",x"48",
x"C9",x"80",x"F0",x"06",x"C9",x"7F",x"F0",x"0D",
x"38",x"24",x"18",x"A9",x"FD",x"20",x"A2",x"F9",
x"A9",x"60",x"20",x"94",x"FA",x"20",x"BA",x"FF",
x"F0",x"FB",x"A0",x"01",x"C9",x"0D",x"F0",x"09",
x"C9",x"1D",x"F0",x"14",x"20",x"95",x"F9",x"D0",
x"EC",x"A5",x"EA",x"91",x"E0",x"20",x"A2",x"FA",
x"A5",x"E3",x"85",x"E0",x"A5",x"E4",x"85",x"E1",
x"A9",x"60",x"85",x"EA",x"91",x"E3",x"E6",x"E3",
x"F0",x"02",x"C6",x"E4",x"88",x"88",x"D1",x"E3",
x"D0",x"FB",x"A2",x"00",x"C8",x"F0",x"0E",x"C0",
x"B6",x"B0",x"02",x"A0",x"B6",x"B1",x"E3",x"95",
x"13",x"E8",x"C8",x"D0",x"F8",x"94",x"13",x"20",
x"BF",x"FA",x"4C",x"6A",x"A8",x"00",x"F0",x"D1",
x"85",x"E2",x"48",x"8A",x"48",x"98",x"48",x"A5",
x"E2",x"A0",x"00",x"84",x"E2",x"20",x"6C",x"FF",
x"C9",x"EC",x"D0",x"1E",x"A9",x"FF",x"2C",x"A9",
x"E0",x"18",x"65",x"E0",x"85",x"E0",x"B0",x"02",
x"C6",x"E1",x"20",x"B1",x"FA",x"A5",x"E0",x"38",
x"E9",x"3F",x"A5",x"E1",x"E9",x"D0",x"90",x"0E",
x"B0",x"44",x"C9",x"1A",x"F0",x"E1",x"C9",x"0A",
x"F0",x"07",x"C9",x"EE",x"D0",x"3A",x"A9",x"01",
x"2C",x"A9",x"20",x"18",x"65",x"E0",x"85",x"E0",
x"90",x"02",x"E6",x"E1",x"20",x"B1",x"FA",x"38",
x"A9",x"9E",x"E5",x"E0",x"A9",x"D3",x"E5",x"E1",
x"B0",x"1C",x"A9",x"60",x"91",x"E0",x"AD",x"22",
x"02",x"F0",x"2D",x"20",x"F1",x"F8",x"30",x"AF",
x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",
x"EA",x"20",x"C8",x"FA",x"90",x"A1",x"A9",x"02",
x"C9",x"0D",x"F0",x"04",x"C9",x"01",x"D0",x"0C",
x"A9",x"1F",x"24",x"E0",x"F0",x"04",x"C6",x"E0",
x"D0",x"F8",x"F0",x"C0",x"C9",x"7F",x"D0",x"0A",
x"A9",x"40",x"A0",x"D0",x"84",x"E1",x"85",x"E0",
x"D0",x"B2",x"C9",x"09",x"D0",x"1C",x"20",x"9C",
x"F9",x"20",x"A0",x"FA",x"C8",x"A5",x"E0",x"85",
x"E5",x"A5",x"E1",x"85",x"E6",x"A5",x"E3",x"A6",
x"E4",x"20",x"DE",x"FA",x"20",x"BB",x"FA",x"B0",
x"85",x"00",x"C9",x"04",x"D0",x"24",x"A0",x"02",
x"B1",x"E0",x"85",x"EA",x"20",x"A0",x"FA",x"A5",
x"E3",x"85",x"E5",x"A5",x"E4",x"85",x"E6",x"A5",
x"E0",x"A6",x"E1",x"69",x"00",x"90",x"01",x"E8",
x"C8",x"20",x"C8",x"FA",x"20",x"BB",x"FA",x"4C",
x"D4",x"F9",x"48",x"A9",x"BF",x"8D",x"00",x"DF",
x"AD",x"00",x"DF",x"29",x"04",x"D0",x"03",x"20",
x"95",x"FC",x"A9",x"FE",x"8D",x"00",x"DF",x"2C",
x"00",x"DF",x"10",x"FB",x"68",x"EA",x"EA",x"EA",
x"EA",x"C9",x"04",x"30",x"0C",x"20",x"99",x"A3",
x"24",x"64",x"30",x"05",x"85",x"EA",x"4C",x"C6",
x"F9",x"A5",x"E2",x"D0",x"08",x"4C",x"6D",x"BF",
x"A0",x"00",x"B1",x"E3",x"C9",x"60",x"F0",x"08",
x"E6",x"E3",x"D0",x"02",x"E6",x"E4",x"D0",x"F2",
x"60",x"A0",x"01",x"A5",x"EA",x"91",x"E3",x"B1",
x"E0",x"85",x"EA",x"A9",x"BB",x"91",x"E0",x"A5",
x"E0",x"85",x"E3",x"A5",x"E1",x"85",x"E4",x"60",
x"85",x"E7",x"86",x"E8",x"A2",x"00",x"B1",x"E7",
x"81",x"E7",x"E6",x"E7",x"D0",x"02",x"E6",x"E8",
x"20",x"F6",x"FA",x"B0",x"F1",x"60",x"85",x"E7",
x"86",x"E8",x"A2",x"00",x"A1",x"E7",x"91",x"E7",
x"A5",x"E7",x"D0",x"02",x"C6",x"E8",x"C6",x"E7",
x"20",x"F6",x"FA",x"90",x"EF",x"60",x"A5",x"E5",
x"38",x"E5",x"E7",x"A5",x"E6",x"E5",x"E8",x"60",
x"68",x"C9",x"30",x"48",x"D0",x"0D",x"86",x"BF",
x"A0",x"01",x"B1",x"C3",x"20",x"81",x"AD",x"B0",
x"0B",x"A6",x"BF",x"E6",x"C3",x"D0",x"02",x"E6",
x"C4",x"4C",x"C2",x"00",x"A5",x"C3",x"D0",x"02",
x"C6",x"C4",x"C6",x"C3",x"A0",x"FF",x"A2",x"00",
x"C8",x"CA",x"BD",x"00",x"FC",x"F0",x"27",x"38",
x"F1",x"C3",x"F0",x"F4",x"C9",x"80",x"F0",x"0C",
x"A0",x"00",x"CA",x"BD",x"01",x"FC",x"10",x"FA",
x"CA",x"CA",x"D0",x"E6",x"20",x"0F",x"A7",x"68",
x"68",x"68",x"68",x"BD",x"FF",x"FB",x"48",x"BD",
x"FE",x"FB",x"48",x"4C",x"13",x"FB",x"A0",x"01",
x"20",x"0F",x"A7",x"4C",x"11",x"FB",x"EA",x"7B",
x"0E",x"FA",x"35",x"EA",x"20",x"D4",x"AF",x"20",
x"BA",x"FF",x"85",x"13",x"A9",x"2C",x"85",x"12",
x"A9",x"00",x"85",x"14",x"A8",x"A2",x"12",x"4C",
x"55",x"A9",x"20",x"D2",x"FB",x"A9",x"5F",x"A0",
x"FB",x"D0",x"07",x"20",x"D2",x"FB",x"A9",x"90",
x"A0",x"FB",x"20",x"FB",x"B5",x"4C",x"BA",x"B7",
x"86",x"65",x"2E",x"E1",x"00",x"FF",x"8D",x"00",
x"F0",x"A9",x"20",x"4C",x"86",x"F9",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"20",x"AE",x"B3",x"20",x"FB",x"AB",x"8A",
x"EA",x"F0",x"0E",x"A2",x"A3",x"A0",x"18",x"C8",
x"D0",x"FD",x"E8",x"D0",x"F8",x"C6",x"AF",x"D0",
x"F2",x"60",x"6C",x"11",x"00",x"20",x"FC",x"B3",
x"8A",x"20",x"C2",x"FB",x"A8",x"A9",x"00",x"6C",
x"08",x"00",x"20",x"F5",x"AB",x"20",x"B0",x"AA",
x"4C",x"BA",x"B7",x"20",x"AD",x"AA",x"20",x"08",
x"B4",x"20",x"32",x"A4",x"38",x"A5",x"AA",x"E9",
x"01",x"A4",x"AB",x"4C",x"21",x"A6",x"20",x"AE",
x"B3",x"86",x"E5",x"20",x"AB",x"B3",x"A5",x"E5",
x"20",x"2B",x"FC",x"A4",x"C1",x"84",x"E2",x"4C",
x"1C",x"FA",x"20",x"AE",x"B3",x"A0",x"FF",x"C8",
x"84",x"C0",x"F0",x"03",x"20",x"AB",x"B3",x"A4",
x"C0",x"96",x"F0",x"C9",x"2C",x"F0",x"F0",x"A4",
x"F1",x"A5",x"F2",x"29",x"03",x"AA",x"BD",x"26",
x"FC",x"A6",x"F0",x"4C",x"00",x"F8",x"00",x"01",
x"81",x"80",x"00",x"29",x"1F",x"85",x"C0",x"8A",
x"49",x"FF",x"6A",x"6A",x"6A",x"A8",x"29",x"03",
x"09",x"D0",x"85",x"C1",x"98",x"6A",x"29",x"E0",
x"05",x"C0",x"85",x"C0",x"EA",x"60",x"20",x"D2",
x"FB",x"A5",x"AC",x"F0",x"30",x"38",x"E9",x"80",
x"F0",x"2B",x"90",x"1A",x"A8",x"C0",x"08",x"90",
x"20",x"A5",x"AE",x"85",x"AD",x"A5",x"AF",x"85",
x"AE",x"A9",x"00",x"85",x"AF",x"98",x"E9",x"08",
x"D0",x"EA",x"A9",x"80",x"85",x"AC",x"4C",x"D5",
x"B4",x"06",x"AF",x"26",x"AE",x"26",x"AD",x"88",
x"98",x"D0",x"F6",x"F0",x"ED",x"60",x"20",x"AE",
x"B3",x"86",x"F4",x"20",x"AB",x"B3",x"86",x"F5",
x"A5",x"F4",x"4C",x"19",x"FB",x"A2",x"A0",x"A0",
x"80",x"A9",x"00",x"F0",x"06",x"A2",x"D4",x"A0",
x"D0",x"A9",x"60",x"84",x"FF",x"A0",x"00",x"84",
x"FE",x"91",x"FE",x"C8",x"D0",x"FB",x"E6",x"FF",
x"E4",x"FF",x"D0",x"F5",x"60",x"B9",x"20",x"D0",
x"99",x"00",x"D0",x"4C",x"01",x"F9",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"28",
x"02",x"C2",x"55",x"53",x"8C",x"FC",x"C7",x"4C",
x"43",x"ED",x"FB",x"D2",x"43",x"53",x"63",x"FB",
x"D4",x"45",x"47",x"94",x"FC",x"C5",x"47",x"41",
x"50",x"A8",x"FB",x"A8",x"59",x"45",x"44",x"DA",
x"FB",x"D4",x"45",x"53",x"82",x"FB",x"C4",x"41",
x"52",x"79",x"FB",x"C7",x"45",x"44",x"45",x"FC",
x"C3",x"41",x"52",x"46",x"C4",x"FB",x"CC",x"4C",
x"41",x"43",x"01",x"FC",x"D3",x"49",x"44",x"47",
x"8A",x"48",x"98",x"48",x"A9",x"01",x"20",x"CD",
x"F8",x"20",x"D5",x"F8",x"D0",x"05",x"0A",x"D0",
x"F5",x"F0",x"53",x"4A",x"90",x"09",x"2A",x"E0",
x"21",x"D0",x"F3",x"A9",x"1B",x"D0",x"21",x"20",
x"C8",x"FD",x"98",x"8D",x"13",x"02",x"0A",x"0A",
x"0A",x"38",x"ED",x"13",x"02",x"8D",x"13",x"02",
x"8A",x"4A",x"20",x"C8",x"FD",x"D0",x"2F",x"18",
x"98",x"6D",x"13",x"02",x"A8",x"B9",x"CF",x"FD",
x"CD",x"15",x"02",x"D0",x"26",x"CE",x"14",x"02",
x"F0",x"2B",x"A0",x"05",x"A2",x"C8",x"CA",x"D0",
x"FD",x"88",x"D0",x"F8",x"F0",x"AE",x"C9",x"01",
x"F0",x"35",x"A0",x"00",x"C9",x"02",x"F0",x"47",
x"A0",x"C0",x"C9",x"20",x"F0",x"41",x"A9",x"00",
x"8D",x"16",x"02",x"8D",x"15",x"02",x"A9",x"02",
x"8D",x"14",x"02",x"D0",x"8F",x"A2",x"96",x"CD",
x"16",x"02",x"D0",x"02",x"A2",x"14",x"8E",x"14",
x"02",x"8D",x"16",x"02",x"A9",x"01",x"20",x"CD",
x"F8",x"20",x"DE",x"F8",x"4A",x"90",x"33",x"AA",
x"29",x"03",x"F0",x"0B",x"A0",x"10",x"AD",x"15",
x"02",x"10",x"0C",x"A0",x"F0",x"D0",x"08",x"A0",
x"00",x"E0",x"20",x"D0",x"02",x"A0",x"C0",x"AD",
x"15",x"02",x"29",x"7F",x"C9",x"20",x"F0",x"07",
x"8C",x"13",x"02",x"18",x"6D",x"13",x"02",x"8D",
x"13",x"02",x"68",x"A8",x"68",x"AA",x"AD",x"13",
x"02",x"60",x"D0",x"92",x"A0",x"20",x"D0",x"DF",
x"A0",x"08",x"88",x"0A",x"90",x"FC",x"60",x"D0",
x"BB",x"2F",x"20",x"5A",x"41",x"51",x"2C",x"4D",
x"4E",x"42",x"56",x"43",x"58",x"4B",x"4A",x"48",
x"47",x"46",x"44",x"53",x"49",x"55",x"59",x"54",
x"52",x"45",x"57",x"00",x"00",x"0D",x"0A",x"4F",
x"4C",x"2E",x"00",x"FF",x"2D",x"BA",x"30",x"B9",
x"B8",x"B7",x"B6",x"B5",x"B4",x"B3",x"B2",x"B1",
x"A2",x"28",x"9A",x"D8",x"A0",x"00",x"A9",x"60",
x"99",x"00",x"D0",x"99",x"00",x"D1",x"99",x"00",
x"D2",x"99",x"00",x"D3",x"C8",x"D0",x"F1",x"F0",
x"19",x"20",x"E9",x"FE",x"C9",x"2F",x"F0",x"1E",
x"C9",x"47",x"F0",x"17",x"C9",x"4C",x"F0",x"59",
x"20",x"93",x"FE",x"30",x"EC",x"A2",x"02",x"20",
x"DA",x"FE",x"B1",x"FE",x"85",x"FC",x"20",x"AC",
x"FE",x"D0",x"DE",x"6C",x"FE",x"00",x"20",x"E9",
x"FE",x"C9",x"2E",x"F0",x"D4",x"C9",x"1D",x"D0",
x"0B",x"A5",x"FE",x"D0",x"02",x"C6",x"FF",x"C6",
x"FE",x"18",x"90",x"11",x"C9",x"0D",x"D0",x"16",
x"A5",x"FB",x"D0",x"03",x"20",x"F1",x"F8",x"E6",
x"FE",x"D0",x"02",x"E6",x"FF",x"A0",x"00",x"B1",
x"FE",x"85",x"FC",x"18",x"90",x"0E",x"20",x"93",
x"FE",x"30",x"CB",x"A2",x"00",x"20",x"DA",x"FE",
x"A5",x"FC",x"91",x"FE",x"20",x"AC",x"FE",x"D0",
x"BD",x"85",x"FB",x"F0",x"B9",x"AD",x"00",x"F0",
x"4A",x"90",x"FA",x"AD",x"01",x"F0",x"29",x"7F",
x"60",x"EA",x"EA",x"C9",x"30",x"30",x"12",x"C9",
x"3A",x"30",x"0B",x"C9",x"41",x"30",x"0A",x"C9",
x"47",x"10",x"06",x"38",x"E9",x"07",x"29",x"0F",
x"60",x"A9",x"80",x"60",x"A2",x"03",x"A0",x"00",
x"B5",x"FC",x"4A",x"4A",x"4A",x"4A",x"20",x"CA",
x"FE",x"B5",x"FC",x"20",x"CA",x"FE",x"CA",x"10",
x"EF",x"A9",x"60",x"8D",x"4A",x"D3",x"8D",x"4B",
x"D3",x"60",x"29",x"0F",x"09",x"30",x"C9",x"3A",
x"30",x"03",x"18",x"69",x"07",x"99",x"46",x"D3",
x"C8",x"60",x"A0",x"04",x"0A",x"0A",x"0A",x"0A",
x"2A",x"36",x"FC",x"36",x"FD",x"88",x"D0",x"F8",
x"60",x"A5",x"FB",x"D0",x"98",x"4C",x"00",x"FD",
x"18",x"F9",x"86",x"F9",x"9B",x"FF",x"8B",x"FF",
x"86",x"F9",x"26",x"02",x"00",x"FE",x"23",x"02",
x"D8",x"A2",x"28",x"9A",x"A0",x"0B",x"B9",x"EF",
x"FE",x"99",x"17",x"02",x"88",x"D0",x"F7",x"8C",
x"06",x"02",x"8C",x"12",x"02",x"8C",x"03",x"02",
x"8C",x"05",x"02",x"20",x"AD",x"F8",x"AD",x"E0",
x"FF",x"8D",x"00",x"02",x"A9",x"60",x"99",x"00",
x"D3",x"99",x"00",x"D2",x"99",x"00",x"D1",x"99",
x"00",x"D0",x"C8",x"D0",x"F1",x"B9",x"5F",x"FF",
x"F0",x"06",x"20",x"86",x"F9",x"C8",x"D0",x"F5",
x"20",x"BA",x"FF",x"C9",x"4D",x"D0",x"03",x"4C",
x"00",x"FE",x"C9",x"57",x"D0",x"03",x"4C",x"00",
x"00",x"C9",x"43",x"D0",x"03",x"4C",x"11",x"BD",
x"C9",x"42",x"D0",x"A4",x"4C",x"E4",x"F8",x"42",
x"2F",x"43",x"2F",x"57",x"2F",x"4D",x"20",x"3F",
x"00",x"20",x"2D",x"BF",x"48",x"AD",x"05",x"02",
x"F0",x"22",x"68",x"20",x"C0",x"F8",x"C9",x"0D",
x"D0",x"1B",x"48",x"8A",x"48",x"A2",x"0A",x"A9",
x"00",x"20",x"C0",x"F8",x"CA",x"D0",x"FA",x"68",
x"AA",x"68",x"60",x"48",x"CE",x"03",x"02",x"A9",
x"00",x"8D",x"05",x"02",x"68",x"60",x"48",x"A9",
x"01",x"D0",x"F6",x"AD",x"12",x"02",x"D0",x"19",
x"A9",x"FE",x"8D",x"00",x"DF",x"2C",x"00",x"DF",
x"70",x"0F",x"A9",x"FB",x"8D",x"00",x"DF",x"2C",
x"00",x"DF",x"70",x"05",x"A9",x"03",x"4C",x"36",
x"A6",x"60",x"2C",x"03",x"02",x"10",x"19",x"A9",
x"FD",x"8D",x"00",x"DF",x"A9",x"10",x"2C",x"00",
x"DF",x"F0",x"0A",x"AD",x"00",x"F0",x"4A",x"90",
x"EE",x"AD",x"01",x"F0",x"60",x"EE",x"03",x"02",
x"4C",x"00",x"FD",x"4C",x"00",x"FB",x"FF",x"FF",
x"60",x"1F",x"00",x"00",x"03",x"FF",x"9F",x"00",
x"03",x"FF",x"9F",x"6C",x"18",x"02",x"6C",x"1A",
x"02",x"6C",x"1C",x"02",x"6C",x"1E",x"02",x"6C",
x"20",x"02",x"26",x"02",x"00",x"FF",x"23",x"02"
);
begin
process (address)
begin
q <= romdata (to_integer(unsigned(address)));
end process;
end behavior;

